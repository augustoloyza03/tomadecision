library verilog;
use verilog.vl_types.all;
entity decision_vlg_vec_tst is
end decision_vlg_vec_tst;
