library verilog;
use verilog.vl_types.all;
entity decisionfinal_vlg_vec_tst is
end decisionfinal_vlg_vec_tst;
